

module collision(enable, x_in, y_in, x_out, y_out, vertical_in, verical_out, horizontal_in, horizontal_out);





endmodule
